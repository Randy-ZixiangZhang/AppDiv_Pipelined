library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.ALL;

entity AppDiv_ROM is
   generic(BIT_WIDTH : integer);
   Port ( clk : in bit;
       addr : in std_logic_vector(8 downto 0);
       data : out unsigned(35 downto 0)
       );
end AppDiv_ROM;

architecture behavioral of AppDiv_ROM is
type rom_type is array (0 to 109) of unsigned(35 downto 0);
signal ROM : rom_type := (
"010000000000001111010000001111010000",
"010000000101001111010000010000101101",
"010000000000001101111011001101111011",
"010000001010001111010000010010001010",
"010000001100001101111011001111001001",
"010000000000001100110011001100110100",
"010000001110001111010000010011100111",
"010000011000001101111011010000010110",
"010000010001001100110011001101110101",
"010000000000001011110110001011110111",
"010000010011001111010000010101000100",
"010000100011001101111011010001100100",
"010000100001001100110011001110110111",
"010000010100001011110110001100101111",
"010000000000001011000010001011000010",
"010000011000001111010000010110100001",
"010000101111001101111011010010110001",
"010000110001001100110011001111111000",
"010000101000001011110110001101100111",
"010000010110001011000010001011110011",
"010000000000001010010100001010010101",
"010000011100001111010000010111111110",
"010000111011001101111011010011111111",
"010001000010001100110011010000111010",
"010000111011001011110110001110011111",
"010000101100001011000010001100100100",
"010000011000001010010100001010111111",
"010000000000001001101100001001101101",
"010000100001001111010000011001011100",
"010001000110001101111011010101001100",
"010001010010001100110011010001111100",
"010001001111001011110110001111011000",
"010001000010001011000010001101010101",
"010000101111001010010100001011101010",
"010000011000001001101100001010010010",
"010000000000001001001001001001001001",
"010000100110001111010000011010111001",
"010001010010001101111011010110011010",
"010001100011001100110011010010111101",
"010001100011001011110110010000010000",
"010001011000001011000010001110000101",
"010001000110001010010100001100010101",
"010000110001001001101100001010111000",
"010000011001001001001001001001101010",
"010000000000001000101001001000101001",
"010000101010001111010000011100010110",
"010001011101001101111011010111100111",
"010001110011001100110011010011111111",
"010001110110001011110110010001001000",
"010001101110001011000010001110110110",
"010001011110001010010100001100111111",
"010001001001001001101100001011011101",
"010000110010001001001001001010001100",
"010000011001001000101001001001000111",
"010000000000001000001101001000001101",
"100000000001011110100000011110100001",
"011111101010011011110110011001011100",
"100000000001011011110110011011110111",
"011110111111011001100111010101100001",
"011111100000011001100111010111100101",
"100000000001011001100111011001101000",
"011110001011010111101101010010011101",
"011110110010010111101101010100001101",
"011111011001010111101101010101111110",
"100000000001010111101101010111101110",
"011101010001010110000101001111111111",
"011101111101010110000101010001100001",
"011110101001010110000101010011000010",
"011111010101010110000101010100100100",
"100000000001010110000101010110000101",
"011100010110010100101001001101111111",
"011101000101010100101001001111010101",
"011101110100010100101001010000101010",
"011110100011010100101001010001111111",
"011111010010010100101001010011010100",
"100000000001010100101001010100101010",
"011011011011010011011001001100010110",
"011100001100010011011001001101100001",
"011100111101010011011001001110101100",
"011101101110010011011001001111111000",
"011110011111010011011001010001000011",
"011111010000010011011001010010001110",
"100000000000010011011001010011011010",
"011010100001010010010010001010111110",
"011011010011010010010010001100000001",
"011100000101010010010010001101000100",
"011100111000010010010010001110000111",
"011101101010010010010010001111001010",
"011110011100010010010010010000001101",
"011111001110010010010010010001010000",
"100000000000010010010010010010010010",
"011001101001010001010011001001110100",
"011010011100010001010011001010110000",
"011011001111010001010011001011101100",
"011100000010010001010011001100101000",
"011100110101010001010011001101100100",
"011101101000010001010011001110011111",
"011110011011010001010011001111011011",
"011111001101010001010011010000010111",
"100000000000010001010011010001010011",
"011000110100010000011010001000110101",
"011001100111010000011010001001101011",
"011010011010010000011010001010100001",
"011011001101010000011010001011010111",
"011100000000010000011010001100001101",
"011100110011010000011010001101000011",
"011101100111010000011010001101111001",
"011110011010010000011010001110101110",
"011111001101010000011010001111100100",
"100000000000010000011010010000011010");
    attribute rom_style : string;
    attribute rom_style of ROM : signal is "block";
begin
   process(clk)
   begin
       if rising_edge(clk) then
           data <= ROM(conv_integer(std_logic_vector(addr)));
       end if;
   end process;
end behavioral;
